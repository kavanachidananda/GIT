module d_tb;
reg clk,reset,d;
wire d;
endmodule

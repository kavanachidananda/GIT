module t_ff(input clk,reset,t,output reg q);

endmodule

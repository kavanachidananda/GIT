module d_tb;

endmodule
